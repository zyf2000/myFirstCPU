/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ROM_ROM                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ROM_ROM( Address,
                Data);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[9:0]  Address;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] Data;
   reg[31:0] Data;

   always @ (Address)
   begin
      case(Address)
         0 : Data = 537985025;
         1 : Data = 134220805;
         2 : Data = 537985025;
         3 : Data = 538050562;
         4 : Data = 538116099;
         5 : Data = 134220809;
         6 : Data = 537985025;
         7 : Data = 538050562;
         8 : Data = 538116099;
         9 : Data = 134220813;
         10 : Data = 537985025;
         11 : Data = 538050562;
         12 : Data = 538116099;
         13 : Data = 134220817;
         14 : Data = 537985025;
         15 : Data = 538050562;
         16 : Data = 538116099;
         17 : Data = 201329929;
         18 : Data = 537919489;
         19 : Data = 537985025;
         20 : Data = 1150912;
         21 : Data = 1122336;
         22 : Data = 537002018;
         23 : Data = 12;
         24 : Data = 1149058;
         25 : Data = 304087041;
         26 : Data = 134220821;
         27 : Data = 1122336;
         28 : Data = 537002018;
         29 : Data = 12;
         30 : Data = 537985025;
         31 : Data = 1149056;
         32 : Data = 1122336;
         33 : Data = 537002018;
         34 : Data = 12;
         35 : Data = 304087041;
         36 : Data = 134220831;
         37 : Data = 537985025;
         38 : Data = 1150912;
         39 : Data = 1122336;
         40 : Data = 537002018;
         41 : Data = 12;
         42 : Data = 1149123;
         43 : Data = 1122336;
         44 : Data = 537002018;
         45 : Data = 12;
         46 : Data = 1149187;
         47 : Data = 1122336;
         48 : Data = 537002018;
         49 : Data = 12;
         50 : Data = 1149187;
         51 : Data = 1122336;
         52 : Data = 537002018;
         53 : Data = 12;
         54 : Data = 1149187;
         55 : Data = 1122336;
         56 : Data = 537002018;
         57 : Data = 12;
         58 : Data = 1149187;
         59 : Data = 1122336;
         60 : Data = 537002018;
         61 : Data = 12;
         62 : Data = 1149187;
         63 : Data = 1122336;
         64 : Data = 537002018;
         65 : Data = 12;
         66 : Data = 1149187;
         67 : Data = 1122336;
         68 : Data = 537002018;
         69 : Data = 12;
         70 : Data = 1149187;
         71 : Data = 1122336;
         72 : Data = 537002018;
         73 : Data = 12;
         74 : Data = 537919489;
         75 : Data = 1089472;
         76 : Data = 1286083;
         77 : Data = 32801;
         78 : Data = 538050572;
         79 : Data = 605421571;
         80 : Data = 638582785;
         81 : Data = 839909391;
         82 : Data = 537395208;
         83 : Data = 537460737;
         84 : Data = 1284352;
         85 : Data = 40933413;
         86 : Data = 1253408;
         87 : Data = 537002018;
         88 : Data = 12;
         89 : Data = 17383458;
         90 : Data = 352387065;
         91 : Data = 571473921;
         92 : Data = 538443791;
         93 : Data = 35160100;
         94 : Data = 1083136;
         95 : Data = 537395208;
         96 : Data = 537460737;
         97 : Data = 1284354;
         98 : Data = 40933413;
         99 : Data = 1253409;
         100 : Data = 537002018;
         101 : Data = 12;
         102 : Data = 17383458;
         103 : Data = 352387065;
         104 : Data = 1083138;
         105 : Data = 46772258;
         106 : Data = 314572801;
         107 : Data = 134220880;
         108 : Data = 16416;
         109 : Data = 17317927;
         110 : Data = 541696;
         111 : Data = 889782271;
         112 : Data = 532513;
         113 : Data = 537002018;
         114 : Data = 12;
         115 : Data = 537985023;
         116 : Data = 537985024;
         117 : Data = -1372585984;
         118 : Data = 571473921;
         119 : Data = 573636612;
         120 : Data = -1372585984;
         121 : Data = 571473921;
         122 : Data = 573636612;
         123 : Data = -1372585984;
         124 : Data = 571473921;
         125 : Data = 573636612;
         126 : Data = -1372585984;
         127 : Data = 571473921;
         128 : Data = 573636612;
         129 : Data = -1372585984;
         130 : Data = 571473921;
         131 : Data = 573636612;
         132 : Data = -1372585984;
         133 : Data = 571473921;
         134 : Data = 573636612;
         135 : Data = -1372585984;
         136 : Data = 571473921;
         137 : Data = 573636612;
         138 : Data = -1372585984;
         139 : Data = 571473921;
         140 : Data = 573636612;
         141 : Data = -1372585984;
         142 : Data = 571473921;
         143 : Data = 573636612;
         144 : Data = -1372585984;
         145 : Data = 571473921;
         146 : Data = 573636612;
         147 : Data = -1372585984;
         148 : Data = 571473921;
         149 : Data = 573636612;
         150 : Data = -1372585984;
         151 : Data = 571473921;
         152 : Data = 573636612;
         153 : Data = -1372585984;
         154 : Data = 571473921;
         155 : Data = 573636612;
         156 : Data = -1372585984;
         157 : Data = 571473921;
         158 : Data = 573636612;
         159 : Data = -1372585984;
         160 : Data = 571473921;
         161 : Data = 573636612;
         162 : Data = -1372585984;
         163 : Data = 571473921;
         164 : Data = 573636612;
         165 : Data = 571473921;
         166 : Data = 32800;
         167 : Data = 537985084;
         168 : Data = -1911357440;
         169 : Data = -1909194752;
         170 : Data = 41173034;
         171 : Data = 285212674;
         172 : Data = -1372389376;
         173 : Data = -1374420992;
         174 : Data = 573702140;
         175 : Data = 370278392;
         176 : Data = 1056800;
         177 : Data = 537002018;
         178 : Data = 12;
         179 : Data = 571473924;
         180 : Data = 537985084;
         181 : Data = 370278386;
         182 : Data = 537002034;
         183 : Data = 12;
         188 : Data = 537395201;
         189 : Data = 537460739;
         190 : Data = 537987190;
         191 : Data = 1150208;
         192 : Data = 1122336;
         193 : Data = 537002018;
         194 : Data = 12;
         195 : Data = 537591816;
         196 : Data = 17926151;
         197 : Data = 20023303;
         198 : Data = 1122336;
         199 : Data = 537002018;
         200 : Data = 12;
         201 : Data = 560726015;
         202 : Data = 358678521;
         203 : Data = 537001994;
         204 : Data = 12;
         209 : Data = 537460735;
         210 : Data = 538015607;
         211 : Data = 1122336;
         212 : Data = 537002018;
         213 : Data = 12;
         214 : Data = 537591824;
         215 : Data = 36210726;
         216 : Data = 1122336;
         217 : Data = 537002018;
         218 : Data = 12;
         219 : Data = 560726015;
         220 : Data = 358678522;
         221 : Data = 537001994;
         222 : Data = 12;
         227 : Data = 537460736;
         228 : Data = 537591824;
         229 : Data = 873563267;
         230 : Data = 538051588;
         231 : Data = 1149952;
         232 : Data = 1217536;
         233 : Data = 909214337;
         234 : Data = 575800324;
         235 : Data = -1389297664;
         236 : Data = 36866080;
         237 : Data = 556335108;
         238 : Data = 560726015;
         239 : Data = 358678523;
         240 : Data = 537591840;
         241 : Data = 537460736;
         242 : Data = -2127495168;
         243 : Data = 1122336;
         244 : Data = 537002018;
         245 : Data = 12;
         246 : Data = 556335105;
         247 : Data = 560726015;
         248 : Data = 358678521;
         249 : Data = 537001994;
         250 : Data = 12;
         255 : Data = 538050545;
         256 : Data = 1122336;
         257 : Data = 537002018;
         258 : Data = 12;
         259 : Data = 573636609;
         260 : Data = 102825979;
         261 : Data = 537001994;
         262 : Data = 12;
         263 : Data = 537001994;
         264 : Data = 12;
         265 : Data = 537919488;
         266 : Data = 571473921;
         267 : Data = 1056800;
         268 : Data = 537002018;
         269 : Data = 12;
         270 : Data = 571473922;
         271 : Data = 1056800;
         272 : Data = 537002018;
         273 : Data = 12;
         274 : Data = 571473923;
         275 : Data = 1056800;
         276 : Data = 537002018;
         277 : Data = 12;
         278 : Data = 571473924;
         279 : Data = 1056800;
         280 : Data = 537002018;
         281 : Data = 12;
         282 : Data = 571473925;
         283 : Data = 1056800;
         284 : Data = 537002018;
         285 : Data = 12;
         286 : Data = 571473926;
         287 : Data = 1056800;
         288 : Data = 537002018;
         289 : Data = 12;
         290 : Data = 571473927;
         291 : Data = 1056800;
         292 : Data = 537002018;
         293 : Data = 12;
         294 : Data = 571473928;
         295 : Data = 1056800;
         296 : Data = 537002018;
         297 : Data = 537002018;
         298 : Data = 12;
         299 : Data = 65011720;
         default : Data = 0;
      endcase
   end

endmodule
